module log_sqrt_lut (
    input wire [15:0] addr,
    output wire signed [7:0] log_sqrt_out  // 2^5 量化
);
    reg signed [7:0] log_sqrt[0:1023];
    initial begin
        log_sqrt[0] = 8'd119;
        log_sqrt[1] = 8'd113;
        log_sqrt[2] = 8'd109;
        log_sqrt[3] = 8'd106;
        log_sqrt[4] = 8'd104;
        log_sqrt[5] = 8'd102;
        log_sqrt[6] = 8'd101;
        log_sqrt[7] = 8'd99;
        log_sqrt[8] = 8'd98;
        log_sqrt[9] = 8'd97;
        log_sqrt[10] = 8'd96;
        log_sqrt[11] = 8'd95;
        log_sqrt[12] = 8'd94;
        log_sqrt[13] = 8'd93;
        log_sqrt[14] = 8'd93;
        log_sqrt[15] = 8'd92;
        log_sqrt[16] = 8'd91;
        log_sqrt[17] = 8'd90;
        log_sqrt[18] = 8'd90;
        log_sqrt[19] = 8'd89;
        log_sqrt[20] = 8'd89;
        log_sqrt[21] = 8'd88;
        log_sqrt[22] = 8'd88;
        log_sqrt[23] = 8'd87;
        log_sqrt[24] = 8'd87;
        log_sqrt[25] = 8'd86;
        log_sqrt[26] = 8'd86;
        log_sqrt[27] = 8'd85;
        log_sqrt[28] = 8'd85;
        log_sqrt[29] = 8'd85;
        log_sqrt[30] = 8'd84;
        log_sqrt[31] = 8'd84;
        log_sqrt[32] = 8'd83;
        log_sqrt[33] = 8'd83;
        log_sqrt[34] = 8'd83;
        log_sqrt[35] = 8'd82;
        log_sqrt[36] = 8'd82;
        log_sqrt[37] = 8'd82;
        log_sqrt[38] = 8'd81;
        log_sqrt[39] = 8'd81;
        log_sqrt[40] = 8'd81;
        log_sqrt[41] = 8'd80;
        log_sqrt[42] = 8'd80;
        log_sqrt[43] = 8'd80;
        log_sqrt[44] = 8'd79;
        log_sqrt[45] = 8'd79;
        log_sqrt[46] = 8'd79;
        log_sqrt[47] = 8'd79;
        log_sqrt[48] = 8'd78;
        log_sqrt[49] = 8'd78;
        log_sqrt[50] = 8'd78;
        log_sqrt[51] = 8'd78;
        log_sqrt[52] = 8'd77;
        log_sqrt[53] = 8'd77;
        log_sqrt[54] = 8'd77;
        log_sqrt[55] = 8'd77;
        log_sqrt[56] = 8'd76;
        log_sqrt[57] = 8'd76;
        log_sqrt[58] = 8'd76;
        log_sqrt[59] = 8'd76;
        log_sqrt[60] = 8'd76;
        log_sqrt[61] = 8'd75;
        log_sqrt[62] = 8'd75;
        log_sqrt[63] = 8'd75;
        log_sqrt[64] = 8'd75;
        log_sqrt[65] = 8'd74;
        log_sqrt[66] = 8'd74;
        log_sqrt[67] = 8'd74;
        log_sqrt[68] = 8'd74;
        log_sqrt[69] = 8'd74;
        log_sqrt[70] = 8'd73;
        log_sqrt[71] = 8'd73;
        log_sqrt[72] = 8'd73;
        log_sqrt[73] = 8'd73;
        log_sqrt[74] = 8'd73;
        log_sqrt[75] = 8'd72;
        log_sqrt[76] = 8'd72;
        log_sqrt[77] = 8'd72;
        log_sqrt[78] = 8'd72;
        log_sqrt[79] = 8'd72;
        log_sqrt[80] = 8'd72;
        log_sqrt[81] = 8'd71;
        log_sqrt[82] = 8'd71;
        log_sqrt[83] = 8'd71;
        log_sqrt[84] = 8'd71;
        log_sqrt[85] = 8'd71;
        log_sqrt[86] = 8'd71;
        log_sqrt[87] = 8'd70;
        log_sqrt[88] = 8'd70;
        log_sqrt[89] = 8'd70;
        log_sqrt[90] = 8'd70;
        log_sqrt[91] = 8'd70;
        log_sqrt[92] = 8'd70;
        log_sqrt[93] = 8'd69;
        log_sqrt[94] = 8'd69;
        log_sqrt[95] = 8'd69;
        log_sqrt[96] = 8'd69;
        log_sqrt[97] = 8'd69;
        log_sqrt[98] = 8'd69;
        log_sqrt[99] = 8'd69;
        log_sqrt[100] = 8'd68;
        log_sqrt[101] = 8'd68;
        log_sqrt[102] = 8'd68;
        log_sqrt[103] = 8'd68;
        log_sqrt[104] = 8'd68;
        log_sqrt[105] = 8'd68;
        log_sqrt[106] = 8'd68;
        log_sqrt[107] = 8'd67;
        log_sqrt[108] = 8'd67;
        log_sqrt[109] = 8'd67;
        log_sqrt[110] = 8'd67;
        log_sqrt[111] = 8'd67;
        log_sqrt[112] = 8'd67;
        log_sqrt[113] = 8'd67;
        log_sqrt[114] = 8'd66;
        log_sqrt[115] = 8'd66;
        log_sqrt[116] = 8'd66;
        log_sqrt[117] = 8'd66;
        log_sqrt[118] = 8'd66;
        log_sqrt[119] = 8'd66;
        log_sqrt[120] = 8'd66;
        log_sqrt[121] = 8'd66;
        log_sqrt[122] = 8'd65;
        log_sqrt[123] = 8'd65;
        log_sqrt[124] = 8'd65;
        log_sqrt[125] = 8'd65;
        log_sqrt[126] = 8'd65;
        log_sqrt[127] = 8'd65;
        log_sqrt[128] = 8'd65;
        log_sqrt[129] = 8'd65;
        log_sqrt[130] = 8'd64;
        log_sqrt[131] = 8'd64;
        log_sqrt[132] = 8'd64;
        log_sqrt[133] = 8'd64;
        log_sqrt[134] = 8'd64;
        log_sqrt[135] = 8'd64;
        log_sqrt[136] = 8'd64;
        log_sqrt[137] = 8'd64;
        log_sqrt[138] = 8'd63;
        log_sqrt[139] = 8'd63;
        log_sqrt[140] = 8'd63;
        log_sqrt[141] = 8'd63;
        log_sqrt[142] = 8'd63;
        log_sqrt[143] = 8'd63;
        log_sqrt[144] = 8'd63;
        log_sqrt[145] = 8'd63;
        log_sqrt[146] = 8'd63;
        log_sqrt[147] = 8'd62;
        log_sqrt[148] = 8'd62;
        log_sqrt[149] = 8'd62;
        log_sqrt[150] = 8'd62;
        log_sqrt[151] = 8'd62;
        log_sqrt[152] = 8'd62;
        log_sqrt[153] = 8'd62;
        log_sqrt[154] = 8'd62;
        log_sqrt[155] = 8'd62;
        log_sqrt[156] = 8'd61;
        log_sqrt[157] = 8'd61;
        log_sqrt[158] = 8'd61;
        log_sqrt[159] = 8'd61;
        log_sqrt[160] = 8'd61;
        log_sqrt[161] = 8'd61;
        log_sqrt[162] = 8'd61;
        log_sqrt[163] = 8'd61;
        log_sqrt[164] = 8'd61;
        log_sqrt[165] = 8'd61;
        log_sqrt[166] = 8'd60;
        log_sqrt[167] = 8'd60;
        log_sqrt[168] = 8'd60;
        log_sqrt[169] = 8'd60;
        log_sqrt[170] = 8'd60;
        log_sqrt[171] = 8'd60;
        log_sqrt[172] = 8'd60;
        log_sqrt[173] = 8'd60;
        log_sqrt[174] = 8'd60;
        log_sqrt[175] = 8'd60;
        log_sqrt[176] = 8'd59;
        log_sqrt[177] = 8'd59;
        log_sqrt[178] = 8'd59;
        log_sqrt[179] = 8'd59;
        log_sqrt[180] = 8'd59;
        log_sqrt[181] = 8'd59;
        log_sqrt[182] = 8'd59;
        log_sqrt[183] = 8'd59;
        log_sqrt[184] = 8'd59;
        log_sqrt[185] = 8'd59;
        log_sqrt[186] = 8'd59;
        log_sqrt[187] = 8'd58;
        log_sqrt[188] = 8'd58;
        log_sqrt[189] = 8'd58;
        log_sqrt[190] = 8'd58;
        log_sqrt[191] = 8'd58;
        log_sqrt[192] = 8'd58;
        log_sqrt[193] = 8'd58;
        log_sqrt[194] = 8'd58;
        log_sqrt[195] = 8'd58;
        log_sqrt[196] = 8'd58;
        log_sqrt[197] = 8'd58;
        log_sqrt[198] = 8'd57;
        log_sqrt[199] = 8'd57;
        log_sqrt[200] = 8'd57;
        log_sqrt[201] = 8'd57;
        log_sqrt[202] = 8'd57;
        log_sqrt[203] = 8'd57;
        log_sqrt[204] = 8'd57;
        log_sqrt[205] = 8'd57;
        log_sqrt[206] = 8'd57;
        log_sqrt[207] = 8'd57;
        log_sqrt[208] = 8'd57;
        log_sqrt[209] = 8'd56;
        log_sqrt[210] = 8'd56;
        log_sqrt[211] = 8'd56;
        log_sqrt[212] = 8'd56;
        log_sqrt[213] = 8'd56;
        log_sqrt[214] = 8'd56;
        log_sqrt[215] = 8'd56;
        log_sqrt[216] = 8'd56;
        log_sqrt[217] = 8'd56;
        log_sqrt[218] = 8'd56;
        log_sqrt[219] = 8'd56;
        log_sqrt[220] = 8'd56;
        log_sqrt[221] = 8'd55;
        log_sqrt[222] = 8'd55;
        log_sqrt[223] = 8'd55;
        log_sqrt[224] = 8'd55;
        log_sqrt[225] = 8'd55;
        log_sqrt[226] = 8'd55;
        log_sqrt[227] = 8'd55;
        log_sqrt[228] = 8'd55;
        log_sqrt[229] = 8'd55;
        log_sqrt[230] = 8'd55;
        log_sqrt[231] = 8'd55;
        log_sqrt[232] = 8'd55;
        log_sqrt[233] = 8'd54;
        log_sqrt[234] = 8'd54;
        log_sqrt[235] = 8'd54;
        log_sqrt[236] = 8'd54;
        log_sqrt[237] = 8'd54;
        log_sqrt[238] = 8'd54;
        log_sqrt[239] = 8'd54;
        log_sqrt[240] = 8'd54;
        log_sqrt[241] = 8'd54;
        log_sqrt[242] = 8'd54;
        log_sqrt[243] = 8'd54;
        log_sqrt[244] = 8'd54;
        log_sqrt[245] = 8'd54;
        log_sqrt[246] = 8'd53;
        log_sqrt[247] = 8'd53;
        log_sqrt[248] = 8'd53;
        log_sqrt[249] = 8'd53;
        log_sqrt[250] = 8'd53;
        log_sqrt[251] = 8'd53;
        log_sqrt[252] = 8'd53;
        log_sqrt[253] = 8'd53;
        log_sqrt[254] = 8'd53;
        log_sqrt[255] = 8'd53;
        log_sqrt[256] = 8'd53;
        log_sqrt[257] = 8'd53;
        log_sqrt[258] = 8'd53;
        log_sqrt[259] = 8'd52;
        log_sqrt[260] = 8'd52;
        log_sqrt[261] = 8'd52;
        log_sqrt[262] = 8'd52;
        log_sqrt[263] = 8'd52;
        log_sqrt[264] = 8'd52;
        log_sqrt[265] = 8'd52;
        log_sqrt[266] = 8'd52;
        log_sqrt[267] = 8'd52;
        log_sqrt[268] = 8'd52;
        log_sqrt[269] = 8'd52;
        log_sqrt[270] = 8'd52;
        log_sqrt[271] = 8'd52;
        log_sqrt[272] = 8'd52;
        log_sqrt[273] = 8'd51;
        log_sqrt[274] = 8'd51;
        log_sqrt[275] = 8'd51;
        log_sqrt[276] = 8'd51;
        log_sqrt[277] = 8'd51;
        log_sqrt[278] = 8'd51;
        log_sqrt[279] = 8'd51;
        log_sqrt[280] = 8'd51;
        log_sqrt[281] = 8'd51;
        log_sqrt[282] = 8'd51;
        log_sqrt[283] = 8'd51;
        log_sqrt[284] = 8'd51;
        log_sqrt[285] = 8'd51;
        log_sqrt[286] = 8'd51;
        log_sqrt[287] = 8'd50;
        log_sqrt[288] = 8'd50;
        log_sqrt[289] = 8'd50;
        log_sqrt[290] = 8'd50;
        log_sqrt[291] = 8'd50;
        log_sqrt[292] = 8'd50;
        log_sqrt[293] = 8'd50;
        log_sqrt[294] = 8'd50;
        log_sqrt[295] = 8'd50;
        log_sqrt[296] = 8'd50;
        log_sqrt[297] = 8'd50;
        log_sqrt[298] = 8'd50;
        log_sqrt[299] = 8'd50;
        log_sqrt[300] = 8'd50;
        log_sqrt[301] = 8'd50;
        log_sqrt[302] = 8'd49;
        log_sqrt[303] = 8'd49;
        log_sqrt[304] = 8'd49;
        log_sqrt[305] = 8'd49;
        log_sqrt[306] = 8'd49;
        log_sqrt[307] = 8'd49;
        log_sqrt[308] = 8'd49;
        log_sqrt[309] = 8'd49;
        log_sqrt[310] = 8'd49;
        log_sqrt[311] = 8'd49;
        log_sqrt[312] = 8'd49;
        log_sqrt[313] = 8'd49;
        log_sqrt[314] = 8'd49;
        log_sqrt[315] = 8'd49;
        log_sqrt[316] = 8'd49;
        log_sqrt[317] = 8'd48;
        log_sqrt[318] = 8'd48;
        log_sqrt[319] = 8'd48;
        log_sqrt[320] = 8'd48;
        log_sqrt[321] = 8'd48;
        log_sqrt[322] = 8'd48;
        log_sqrt[323] = 8'd48;
        log_sqrt[324] = 8'd48;
        log_sqrt[325] = 8'd48;
        log_sqrt[326] = 8'd48;
        log_sqrt[327] = 8'd48;
        log_sqrt[328] = 8'd48;
        log_sqrt[329] = 8'd48;
        log_sqrt[330] = 8'd48;
        log_sqrt[331] = 8'd48;
        log_sqrt[332] = 8'd47;
        log_sqrt[333] = 8'd47;
        log_sqrt[334] = 8'd47;
        log_sqrt[335] = 8'd47;
        log_sqrt[336] = 8'd47;
        log_sqrt[337] = 8'd47;
        log_sqrt[338] = 8'd47;
        log_sqrt[339] = 8'd47;
        log_sqrt[340] = 8'd47;
        log_sqrt[341] = 8'd47;
        log_sqrt[342] = 8'd47;
        log_sqrt[343] = 8'd47;
        log_sqrt[344] = 8'd47;
        log_sqrt[345] = 8'd47;
        log_sqrt[346] = 8'd47;
        log_sqrt[347] = 8'd47;
        log_sqrt[348] = 8'd46;
        log_sqrt[349] = 8'd46;
        log_sqrt[350] = 8'd46;
        log_sqrt[351] = 8'd46;
        log_sqrt[352] = 8'd46;
        log_sqrt[353] = 8'd46;
        log_sqrt[354] = 8'd46;
        log_sqrt[355] = 8'd46;
        log_sqrt[356] = 8'd46;
        log_sqrt[357] = 8'd46;
        log_sqrt[358] = 8'd46;
        log_sqrt[359] = 8'd46;
        log_sqrt[360] = 8'd46;
        log_sqrt[361] = 8'd46;
        log_sqrt[362] = 8'd46;
        log_sqrt[363] = 8'd46;
        log_sqrt[364] = 8'd45;
        log_sqrt[365] = 8'd45;
        log_sqrt[366] = 8'd45;
        log_sqrt[367] = 8'd45;
        log_sqrt[368] = 8'd45;
        log_sqrt[369] = 8'd45;
        log_sqrt[370] = 8'd45;
        log_sqrt[371] = 8'd45;
        log_sqrt[372] = 8'd45;
        log_sqrt[373] = 8'd45;
        log_sqrt[374] = 8'd45;
        log_sqrt[375] = 8'd45;
        log_sqrt[376] = 8'd45;
        log_sqrt[377] = 8'd45;
        log_sqrt[378] = 8'd45;
        log_sqrt[379] = 8'd45;
        log_sqrt[380] = 8'd44;
        log_sqrt[381] = 8'd44;
        log_sqrt[382] = 8'd44;
        log_sqrt[383] = 8'd44;
        log_sqrt[384] = 8'd44;
        log_sqrt[385] = 8'd44;
        log_sqrt[386] = 8'd44;
        log_sqrt[387] = 8'd44;
        log_sqrt[388] = 8'd44;
        log_sqrt[389] = 8'd44;
        log_sqrt[390] = 8'd44;
        log_sqrt[391] = 8'd44;
        log_sqrt[392] = 8'd44;
        log_sqrt[393] = 8'd44;
        log_sqrt[394] = 8'd44;
        log_sqrt[395] = 8'd44;
        log_sqrt[396] = 8'd44;
        log_sqrt[397] = 8'd43;
        log_sqrt[398] = 8'd43;
        log_sqrt[399] = 8'd43;
        log_sqrt[400] = 8'd43;
        log_sqrt[401] = 8'd43;
        log_sqrt[402] = 8'd43;
        log_sqrt[403] = 8'd43;
        log_sqrt[404] = 8'd43;
        log_sqrt[405] = 8'd43;
        log_sqrt[406] = 8'd43;
        log_sqrt[407] = 8'd43;
        log_sqrt[408] = 8'd43;
        log_sqrt[409] = 8'd43;
        log_sqrt[410] = 8'd43;
        log_sqrt[411] = 8'd43;
        log_sqrt[412] = 8'd43;
        log_sqrt[413] = 8'd43;
        log_sqrt[414] = 8'd43;
        log_sqrt[415] = 8'd42;
        log_sqrt[416] = 8'd42;
        log_sqrt[417] = 8'd42;
        log_sqrt[418] = 8'd42;
        log_sqrt[419] = 8'd42;
        log_sqrt[420] = 8'd42;
        log_sqrt[421] = 8'd42;
        log_sqrt[422] = 8'd42;
        log_sqrt[423] = 8'd42;
        log_sqrt[424] = 8'd42;
        log_sqrt[425] = 8'd42;
        log_sqrt[426] = 8'd42;
        log_sqrt[427] = 8'd42;
        log_sqrt[428] = 8'd42;
        log_sqrt[429] = 8'd42;
        log_sqrt[430] = 8'd42;
        log_sqrt[431] = 8'd42;
        log_sqrt[432] = 8'd41;
        log_sqrt[433] = 8'd41;
        log_sqrt[434] = 8'd41;
        log_sqrt[435] = 8'd41;
        log_sqrt[436] = 8'd41;
        log_sqrt[437] = 8'd41;
        log_sqrt[438] = 8'd41;
        log_sqrt[439] = 8'd41;
        log_sqrt[440] = 8'd41;
        log_sqrt[441] = 8'd41;
        log_sqrt[442] = 8'd41;
        log_sqrt[443] = 8'd41;
        log_sqrt[444] = 8'd41;
        log_sqrt[445] = 8'd41;
        log_sqrt[446] = 8'd41;
        log_sqrt[447] = 8'd41;
        log_sqrt[448] = 8'd41;
        log_sqrt[449] = 8'd41;
        log_sqrt[450] = 8'd40;
        log_sqrt[451] = 8'd40;
        log_sqrt[452] = 8'd40;
        log_sqrt[453] = 8'd40;
        log_sqrt[454] = 8'd40;
        log_sqrt[455] = 8'd40;
        log_sqrt[456] = 8'd40;
        log_sqrt[457] = 8'd40;
        log_sqrt[458] = 8'd40;
        log_sqrt[459] = 8'd40;
        log_sqrt[460] = 8'd40;
        log_sqrt[461] = 8'd40;
        log_sqrt[462] = 8'd40;
        log_sqrt[463] = 8'd40;
        log_sqrt[464] = 8'd40;
        log_sqrt[465] = 8'd40;
        log_sqrt[466] = 8'd40;
        log_sqrt[467] = 8'd40;
        log_sqrt[468] = 8'd39;
        log_sqrt[469] = 8'd39;
        log_sqrt[470] = 8'd39;
        log_sqrt[471] = 8'd39;
        log_sqrt[472] = 8'd39;
        log_sqrt[473] = 8'd39;
        log_sqrt[474] = 8'd39;
        log_sqrt[475] = 8'd39;
        log_sqrt[476] = 8'd39;
        log_sqrt[477] = 8'd39;
        log_sqrt[478] = 8'd39;
        log_sqrt[479] = 8'd39;
        log_sqrt[480] = 8'd39;
        log_sqrt[481] = 8'd39;
        log_sqrt[482] = 8'd39;
        log_sqrt[483] = 8'd39;
        log_sqrt[484] = 8'd39;
        log_sqrt[485] = 8'd39;
        log_sqrt[486] = 8'd39;
        log_sqrt[487] = 8'd38;
        log_sqrt[488] = 8'd38;
        log_sqrt[489] = 8'd38;
        log_sqrt[490] = 8'd38;
        log_sqrt[491] = 8'd38;
        log_sqrt[492] = 8'd38;
        log_sqrt[493] = 8'd38;
        log_sqrt[494] = 8'd38;
        log_sqrt[495] = 8'd38;
        log_sqrt[496] = 8'd38;
        log_sqrt[497] = 8'd38;
        log_sqrt[498] = 8'd38;
        log_sqrt[499] = 8'd38;
        log_sqrt[500] = 8'd38;
        log_sqrt[501] = 8'd38;
        log_sqrt[502] = 8'd38;
        log_sqrt[503] = 8'd38;
        log_sqrt[504] = 8'd38;
        log_sqrt[505] = 8'd37;
        log_sqrt[506] = 8'd37;
        log_sqrt[507] = 8'd37;
        log_sqrt[508] = 8'd37;
        log_sqrt[509] = 8'd37;
        log_sqrt[510] = 8'd37;
        log_sqrt[511] = 8'd37;
        log_sqrt[512] = 8'd37;
        log_sqrt[513] = 8'd37;
        log_sqrt[514] = 8'd37;
        log_sqrt[515] = 8'd37;
        log_sqrt[516] = 8'd37;
        log_sqrt[517] = 8'd37;
        log_sqrt[518] = 8'd37;
        log_sqrt[519] = 8'd37;
        log_sqrt[520] = 8'd37;
        log_sqrt[521] = 8'd37;
        log_sqrt[522] = 8'd37;
        log_sqrt[523] = 8'd37;
        log_sqrt[524] = 8'd36;
        log_sqrt[525] = 8'd36;
        log_sqrt[526] = 8'd36;
        log_sqrt[527] = 8'd36;
        log_sqrt[528] = 8'd36;
        log_sqrt[529] = 8'd36;
        log_sqrt[530] = 8'd36;
        log_sqrt[531] = 8'd36;
        log_sqrt[532] = 8'd36;
        log_sqrt[533] = 8'd36;
        log_sqrt[534] = 8'd36;
        log_sqrt[535] = 8'd36;
        log_sqrt[536] = 8'd36;
        log_sqrt[537] = 8'd36;
        log_sqrt[538] = 8'd36;
        log_sqrt[539] = 8'd36;
        log_sqrt[540] = 8'd36;
        log_sqrt[541] = 8'd36;
        log_sqrt[542] = 8'd36;
        log_sqrt[543] = 8'd35;
        log_sqrt[544] = 8'd35;
        log_sqrt[545] = 8'd35;
        log_sqrt[546] = 8'd35;
        log_sqrt[547] = 8'd35;
        log_sqrt[548] = 8'd35;
        log_sqrt[549] = 8'd35;
        log_sqrt[550] = 8'd35;
        log_sqrt[551] = 8'd35;
        log_sqrt[552] = 8'd35;
        log_sqrt[553] = 8'd35;
        log_sqrt[554] = 8'd35;
        log_sqrt[555] = 8'd35;
        log_sqrt[556] = 8'd35;
        log_sqrt[557] = 8'd35;
        log_sqrt[558] = 8'd35;
        log_sqrt[559] = 8'd35;
        log_sqrt[560] = 8'd35;
        log_sqrt[561] = 8'd35;
        log_sqrt[562] = 8'd35;
        log_sqrt[563] = 8'd34;
        log_sqrt[564] = 8'd34;
        log_sqrt[565] = 8'd34;
        log_sqrt[566] = 8'd34;
        log_sqrt[567] = 8'd34;
        log_sqrt[568] = 8'd34;
        log_sqrt[569] = 8'd34;
        log_sqrt[570] = 8'd34;
        log_sqrt[571] = 8'd34;
        log_sqrt[572] = 8'd34;
        log_sqrt[573] = 8'd34;
        log_sqrt[574] = 8'd34;
        log_sqrt[575] = 8'd34;
        log_sqrt[576] = 8'd34;
        log_sqrt[577] = 8'd34;
        log_sqrt[578] = 8'd34;
        log_sqrt[579] = 8'd34;
        log_sqrt[580] = 8'd34;
        log_sqrt[581] = 8'd34;
        log_sqrt[582] = 8'd33;
        log_sqrt[583] = 8'd33;
        log_sqrt[584] = 8'd33;
        log_sqrt[585] = 8'd33;
        log_sqrt[586] = 8'd33;
        log_sqrt[587] = 8'd33;
        log_sqrt[588] = 8'd33;
        log_sqrt[589] = 8'd33;
        log_sqrt[590] = 8'd33;
        log_sqrt[591] = 8'd33;
        log_sqrt[592] = 8'd33;
        log_sqrt[593] = 8'd33;
        log_sqrt[594] = 8'd33;
        log_sqrt[595] = 8'd33;
        log_sqrt[596] = 8'd33;
        log_sqrt[597] = 8'd33;
        log_sqrt[598] = 8'd33;
        log_sqrt[599] = 8'd33;
        log_sqrt[600] = 8'd33;
        log_sqrt[601] = 8'd32;
        log_sqrt[602] = 8'd32;
        log_sqrt[603] = 8'd32;
        log_sqrt[604] = 8'd32;
        log_sqrt[605] = 8'd32;
        log_sqrt[606] = 8'd32;
        log_sqrt[607] = 8'd32;
        log_sqrt[608] = 8'd32;
        log_sqrt[609] = 8'd32;
        log_sqrt[610] = 8'd32;
        log_sqrt[611] = 8'd32;
        log_sqrt[612] = 8'd32;
        log_sqrt[613] = 8'd32;
        log_sqrt[614] = 8'd32;
        log_sqrt[615] = 8'd32;
        log_sqrt[616] = 8'd32;
        log_sqrt[617] = 8'd32;
        log_sqrt[618] = 8'd32;
        log_sqrt[619] = 8'd32;
        log_sqrt[620] = 8'd32;
        log_sqrt[621] = 8'd31;
        log_sqrt[622] = 8'd31;
        log_sqrt[623] = 8'd31;
        log_sqrt[624] = 8'd31;
        log_sqrt[625] = 8'd31;
        log_sqrt[626] = 8'd31;
        log_sqrt[627] = 8'd31;
        log_sqrt[628] = 8'd31;
        log_sqrt[629] = 8'd31;
        log_sqrt[630] = 8'd31;
        log_sqrt[631] = 8'd31;
        log_sqrt[632] = 8'd31;
        log_sqrt[633] = 8'd31;
        log_sqrt[634] = 8'd31;
        log_sqrt[635] = 8'd31;
        log_sqrt[636] = 8'd31;
        log_sqrt[637] = 8'd31;
        log_sqrt[638] = 8'd31;
        log_sqrt[639] = 8'd31;
        log_sqrt[640] = 8'd30;
        log_sqrt[641] = 8'd30;
        log_sqrt[642] = 8'd30;
        log_sqrt[643] = 8'd30;
        log_sqrt[644] = 8'd30;
        log_sqrt[645] = 8'd30;
        log_sqrt[646] = 8'd30;
        log_sqrt[647] = 8'd30;
        log_sqrt[648] = 8'd30;
        log_sqrt[649] = 8'd30;
        log_sqrt[650] = 8'd30;
        log_sqrt[651] = 8'd30;
        log_sqrt[652] = 8'd30;
        log_sqrt[653] = 8'd30;
        log_sqrt[654] = 8'd30;
        log_sqrt[655] = 8'd30;
        log_sqrt[656] = 8'd30;
        log_sqrt[657] = 8'd30;
        log_sqrt[658] = 8'd30;
        log_sqrt[659] = 8'd29;
        log_sqrt[660] = 8'd29;
        log_sqrt[661] = 8'd29;
        log_sqrt[662] = 8'd29;
        log_sqrt[663] = 8'd29;
        log_sqrt[664] = 8'd29;
        log_sqrt[665] = 8'd29;
        log_sqrt[666] = 8'd29;
        log_sqrt[667] = 8'd29;
        log_sqrt[668] = 8'd29;
        log_sqrt[669] = 8'd29;
        log_sqrt[670] = 8'd29;
        log_sqrt[671] = 8'd29;
        log_sqrt[672] = 8'd29;
        log_sqrt[673] = 8'd29;
        log_sqrt[674] = 8'd29;
        log_sqrt[675] = 8'd29;
        log_sqrt[676] = 8'd29;
        log_sqrt[677] = 8'd29;
        log_sqrt[678] = 8'd29;
        log_sqrt[679] = 8'd28;
        log_sqrt[680] = 8'd28;
        log_sqrt[681] = 8'd28;
        log_sqrt[682] = 8'd28;
        log_sqrt[683] = 8'd28;
        log_sqrt[684] = 8'd28;
        log_sqrt[685] = 8'd28;
        log_sqrt[686] = 8'd28;
        log_sqrt[687] = 8'd28;
        log_sqrt[688] = 8'd28;
        log_sqrt[689] = 8'd28;
        log_sqrt[690] = 8'd28;
        log_sqrt[691] = 8'd28;
        log_sqrt[692] = 8'd28;
        log_sqrt[693] = 8'd28;
        log_sqrt[694] = 8'd28;
        log_sqrt[695] = 8'd28;
        log_sqrt[696] = 8'd28;
        log_sqrt[697] = 8'd28;
        log_sqrt[698] = 8'd27;
        log_sqrt[699] = 8'd27;
        log_sqrt[700] = 8'd27;
        log_sqrt[701] = 8'd27;
        log_sqrt[702] = 8'd27;
        log_sqrt[703] = 8'd27;
        log_sqrt[704] = 8'd27;
        log_sqrt[705] = 8'd27;
        log_sqrt[706] = 8'd27;
        log_sqrt[707] = 8'd27;
        log_sqrt[708] = 8'd27;
        log_sqrt[709] = 8'd27;
        log_sqrt[710] = 8'd27;
        log_sqrt[711] = 8'd27;
        log_sqrt[712] = 8'd27;
        log_sqrt[713] = 8'd27;
        log_sqrt[714] = 8'd27;
        log_sqrt[715] = 8'd27;
        log_sqrt[716] = 8'd27;
        log_sqrt[717] = 8'd26;
        log_sqrt[718] = 8'd26;
        log_sqrt[719] = 8'd26;
        log_sqrt[720] = 8'd26;
        log_sqrt[721] = 8'd26;
        log_sqrt[722] = 8'd26;
        log_sqrt[723] = 8'd26;
        log_sqrt[724] = 8'd26;
        log_sqrt[725] = 8'd26;
        log_sqrt[726] = 8'd26;
        log_sqrt[727] = 8'd26;
        log_sqrt[728] = 8'd26;
        log_sqrt[729] = 8'd26;
        log_sqrt[730] = 8'd26;
        log_sqrt[731] = 8'd26;
        log_sqrt[732] = 8'd26;
        log_sqrt[733] = 8'd26;
        log_sqrt[734] = 8'd26;
        log_sqrt[735] = 8'd26;
        log_sqrt[736] = 8'd25;
        log_sqrt[737] = 8'd25;
        log_sqrt[738] = 8'd25;
        log_sqrt[739] = 8'd25;
        log_sqrt[740] = 8'd25;
        log_sqrt[741] = 8'd25;
        log_sqrt[742] = 8'd25;
        log_sqrt[743] = 8'd25;
        log_sqrt[744] = 8'd25;
        log_sqrt[745] = 8'd25;
        log_sqrt[746] = 8'd25;
        log_sqrt[747] = 8'd25;
        log_sqrt[748] = 8'd25;
        log_sqrt[749] = 8'd25;
        log_sqrt[750] = 8'd25;
        log_sqrt[751] = 8'd25;
        log_sqrt[752] = 8'd25;
        log_sqrt[753] = 8'd25;
        log_sqrt[754] = 8'd24;
        log_sqrt[755] = 8'd24;
        log_sqrt[756] = 8'd24;
        log_sqrt[757] = 8'd24;
        log_sqrt[758] = 8'd24;
        log_sqrt[759] = 8'd24;
        log_sqrt[760] = 8'd24;
        log_sqrt[761] = 8'd24;
        log_sqrt[762] = 8'd24;
        log_sqrt[763] = 8'd24;
        log_sqrt[764] = 8'd24;
        log_sqrt[765] = 8'd24;
        log_sqrt[766] = 8'd24;
        log_sqrt[767] = 8'd24;
        log_sqrt[768] = 8'd24;
        log_sqrt[769] = 8'd24;
        log_sqrt[770] = 8'd24;
        log_sqrt[771] = 8'd24;
        log_sqrt[772] = 8'd23;
        log_sqrt[773] = 8'd23;
        log_sqrt[774] = 8'd23;
        log_sqrt[775] = 8'd23;
        log_sqrt[776] = 8'd23;
        log_sqrt[777] = 8'd23;
        log_sqrt[778] = 8'd23;
        log_sqrt[779] = 8'd23;
        log_sqrt[780] = 8'd23;
        log_sqrt[781] = 8'd23;
        log_sqrt[782] = 8'd23;
        log_sqrt[783] = 8'd23;
        log_sqrt[784] = 8'd23;
        log_sqrt[785] = 8'd23;
        log_sqrt[786] = 8'd23;
        log_sqrt[787] = 8'd23;
        log_sqrt[788] = 8'd23;
        log_sqrt[789] = 8'd23;
        log_sqrt[790] = 8'd22;
        log_sqrt[791] = 8'd22;
        log_sqrt[792] = 8'd22;
        log_sqrt[793] = 8'd22;
        log_sqrt[794] = 8'd22;
        log_sqrt[795] = 8'd22;
        log_sqrt[796] = 8'd22;
        log_sqrt[797] = 8'd22;
        log_sqrt[798] = 8'd22;
        log_sqrt[799] = 8'd22;
        log_sqrt[800] = 8'd22;
        log_sqrt[801] = 8'd22;
        log_sqrt[802] = 8'd22;
        log_sqrt[803] = 8'd22;
        log_sqrt[804] = 8'd22;
        log_sqrt[805] = 8'd22;
        log_sqrt[806] = 8'd22;
        log_sqrt[807] = 8'd22;
        log_sqrt[808] = 8'd21;
        log_sqrt[809] = 8'd21;
        log_sqrt[810] = 8'd21;
        log_sqrt[811] = 8'd21;
        log_sqrt[812] = 8'd21;
        log_sqrt[813] = 8'd21;
        log_sqrt[814] = 8'd21;
        log_sqrt[815] = 8'd21;
        log_sqrt[816] = 8'd21;
        log_sqrt[817] = 8'd21;
        log_sqrt[818] = 8'd21;
        log_sqrt[819] = 8'd21;
        log_sqrt[820] = 8'd21;
        log_sqrt[821] = 8'd21;
        log_sqrt[822] = 8'd21;
        log_sqrt[823] = 8'd21;
        log_sqrt[824] = 8'd21;
        log_sqrt[825] = 8'd20;
        log_sqrt[826] = 8'd20;
        log_sqrt[827] = 8'd20;
        log_sqrt[828] = 8'd20;
        log_sqrt[829] = 8'd20;
        log_sqrt[830] = 8'd20;
        log_sqrt[831] = 8'd20;
        log_sqrt[832] = 8'd20;
        log_sqrt[833] = 8'd20;
        log_sqrt[834] = 8'd20;
        log_sqrt[835] = 8'd20;
        log_sqrt[836] = 8'd20;
        log_sqrt[837] = 8'd20;
        log_sqrt[838] = 8'd20;
        log_sqrt[839] = 8'd20;
        log_sqrt[840] = 8'd20;
        log_sqrt[841] = 8'd20;
        log_sqrt[842] = 8'd19;
        log_sqrt[843] = 8'd19;
        log_sqrt[844] = 8'd19;
        log_sqrt[845] = 8'd19;
        log_sqrt[846] = 8'd19;
        log_sqrt[847] = 8'd19;
        log_sqrt[848] = 8'd19;
        log_sqrt[849] = 8'd19;
        log_sqrt[850] = 8'd19;
        log_sqrt[851] = 8'd19;
        log_sqrt[852] = 8'd19;
        log_sqrt[853] = 8'd19;
        log_sqrt[854] = 8'd19;
        log_sqrt[855] = 8'd19;
        log_sqrt[856] = 8'd19;
        log_sqrt[857] = 8'd19;
        log_sqrt[858] = 8'd18;
        log_sqrt[859] = 8'd18;
        log_sqrt[860] = 8'd18;
        log_sqrt[861] = 8'd18;
        log_sqrt[862] = 8'd18;
        log_sqrt[863] = 8'd18;
        log_sqrt[864] = 8'd18;
        log_sqrt[865] = 8'd18;
        log_sqrt[866] = 8'd18;
        log_sqrt[867] = 8'd18;
        log_sqrt[868] = 8'd18;
        log_sqrt[869] = 8'd18;
        log_sqrt[870] = 8'd18;
        log_sqrt[871] = 8'd18;
        log_sqrt[872] = 8'd18;
        log_sqrt[873] = 8'd18;
        log_sqrt[874] = 8'd17;
        log_sqrt[875] = 8'd17;
        log_sqrt[876] = 8'd17;
        log_sqrt[877] = 8'd17;
        log_sqrt[878] = 8'd17;
        log_sqrt[879] = 8'd17;
        log_sqrt[880] = 8'd17;
        log_sqrt[881] = 8'd17;
        log_sqrt[882] = 8'd17;
        log_sqrt[883] = 8'd17;
        log_sqrt[884] = 8'd17;
        log_sqrt[885] = 8'd17;
        log_sqrt[886] = 8'd17;
        log_sqrt[887] = 8'd17;
        log_sqrt[888] = 8'd17;
        log_sqrt[889] = 8'd16;
        log_sqrt[890] = 8'd16;
        log_sqrt[891] = 8'd16;
        log_sqrt[892] = 8'd16;
        log_sqrt[893] = 8'd16;
        log_sqrt[894] = 8'd16;
        log_sqrt[895] = 8'd16;
        log_sqrt[896] = 8'd16;
        log_sqrt[897] = 8'd16;
        log_sqrt[898] = 8'd16;
        log_sqrt[899] = 8'd16;
        log_sqrt[900] = 8'd16;
        log_sqrt[901] = 8'd16;
        log_sqrt[902] = 8'd16;
        log_sqrt[903] = 8'd15;
        log_sqrt[904] = 8'd15;
        log_sqrt[905] = 8'd15;
        log_sqrt[906] = 8'd15;
        log_sqrt[907] = 8'd15;
        log_sqrt[908] = 8'd15;
        log_sqrt[909] = 8'd15;
        log_sqrt[910] = 8'd15;
        log_sqrt[911] = 8'd15;
        log_sqrt[912] = 8'd15;
        log_sqrt[913] = 8'd15;
        log_sqrt[914] = 8'd15;
        log_sqrt[915] = 8'd15;
        log_sqrt[916] = 8'd15;
        log_sqrt[917] = 8'd14;
        log_sqrt[918] = 8'd14;
        log_sqrt[919] = 8'd14;
        log_sqrt[920] = 8'd14;
        log_sqrt[921] = 8'd14;
        log_sqrt[922] = 8'd14;
        log_sqrt[923] = 8'd14;
        log_sqrt[924] = 8'd14;
        log_sqrt[925] = 8'd14;
        log_sqrt[926] = 8'd14;
        log_sqrt[927] = 8'd14;
        log_sqrt[928] = 8'd14;
        log_sqrt[929] = 8'd14;
        log_sqrt[930] = 8'd13;
        log_sqrt[931] = 8'd13;
        log_sqrt[932] = 8'd13;
        log_sqrt[933] = 8'd13;
        log_sqrt[934] = 8'd13;
        log_sqrt[935] = 8'd13;
        log_sqrt[936] = 8'd13;
        log_sqrt[937] = 8'd13;
        log_sqrt[938] = 8'd13;
        log_sqrt[939] = 8'd13;
        log_sqrt[940] = 8'd13;
        log_sqrt[941] = 8'd13;
        log_sqrt[942] = 8'd12;
        log_sqrt[943] = 8'd12;
        log_sqrt[944] = 8'd12;
        log_sqrt[945] = 8'd12;
        log_sqrt[946] = 8'd12;
        log_sqrt[947] = 8'd12;
        log_sqrt[948] = 8'd12;
        log_sqrt[949] = 8'd12;
        log_sqrt[950] = 8'd12;
        log_sqrt[951] = 8'd12;
        log_sqrt[952] = 8'd12;
        log_sqrt[953] = 8'd12;
        log_sqrt[954] = 8'd11;
        log_sqrt[955] = 8'd11;
        log_sqrt[956] = 8'd11;
        log_sqrt[957] = 8'd11;
        log_sqrt[958] = 8'd11;
        log_sqrt[959] = 8'd11;
        log_sqrt[960] = 8'd11;
        log_sqrt[961] = 8'd11;
        log_sqrt[962] = 8'd11;
        log_sqrt[963] = 8'd11;
        log_sqrt[964] = 8'd11;
        log_sqrt[965] = 8'd10;
        log_sqrt[966] = 8'd10;
        log_sqrt[967] = 8'd10;
        log_sqrt[968] = 8'd10;
        log_sqrt[969] = 8'd10;
        log_sqrt[970] = 8'd10;
        log_sqrt[971] = 8'd10;
        log_sqrt[972] = 8'd10;
        log_sqrt[973] = 8'd10;
        log_sqrt[974] = 8'd10;
        log_sqrt[975] = 8'd9;
        log_sqrt[976] = 8'd9;
        log_sqrt[977] = 8'd9;
        log_sqrt[978] = 8'd9;
        log_sqrt[979] = 8'd9;
        log_sqrt[980] = 8'd9;
        log_sqrt[981] = 8'd9;
        log_sqrt[982] = 8'd9;
        log_sqrt[983] = 8'd9;
        log_sqrt[984] = 8'd8;
        log_sqrt[985] = 8'd8;
        log_sqrt[986] = 8'd8;
        log_sqrt[987] = 8'd8;
        log_sqrt[988] = 8'd8;
        log_sqrt[989] = 8'd8;
        log_sqrt[990] = 8'd8;
        log_sqrt[991] = 8'd8;
        log_sqrt[992] = 8'd7;
        log_sqrt[993] = 8'd7;
        log_sqrt[994] = 8'd7;
        log_sqrt[995] = 8'd7;
        log_sqrt[996] = 8'd7;
        log_sqrt[997] = 8'd7;
        log_sqrt[998] = 8'd7;
        log_sqrt[999] = 8'd6;
        log_sqrt[1000] = 8'd6;
        log_sqrt[1001] = 8'd6;
        log_sqrt[1002] = 8'd6;
        log_sqrt[1003] = 8'd6;
        log_sqrt[1004] = 8'd6;
        log_sqrt[1005] = 8'd6;
        log_sqrt[1006] = 8'd5;
        log_sqrt[1007] = 8'd5;
        log_sqrt[1008] = 8'd5;
        log_sqrt[1009] = 8'd5;
        log_sqrt[1010] = 8'd5;
        log_sqrt[1011] = 8'd4;
        log_sqrt[1012] = 8'd4;
        log_sqrt[1013] = 8'd4;
        log_sqrt[1014] = 8'd4;
        log_sqrt[1015] = 8'd4;
        log_sqrt[1016] = 8'd3;
        log_sqrt[1017] = 8'd3;
        log_sqrt[1018] = 8'd3;
        log_sqrt[1019] = 8'd2;
        log_sqrt[1020] = 8'd2;
        log_sqrt[1021] = 8'd2;
        log_sqrt[1022] = 8'd1;
        log_sqrt[1023] = 8'd0;
    end
    
    assign log_sqrt_out = log_sqrt[addr[9:0]];

endmodule