module random_gaussian_normal_lut (
    input wire [15:0] addr1,
    input wire [15:0] addr2,
    output wire signed [15:0] random_gaussian_normal_o1,
    output wire signed [15:0] random_gaussian_normal_o2
);
    reg [15:0] random_gaussian_normal[0:1023];
    initial begin
        random_gaussian_normal[0] = 16'd127;
        random_gaussian_normal[1] = 16'd226;
        random_gaussian_normal[2] = 16'd196;
        random_gaussian_normal[3] = 16'd45;
        random_gaussian_normal[4] = 16'd110;
        random_gaussian_normal[5] = 16'd382;
        random_gaussian_normal[6] = 16'd45;
        random_gaussian_normal[7] = 16'd233;
        random_gaussian_normal[8] = 16'd28;
        random_gaussian_normal[9] = 16'd125;
        random_gaussian_normal[10] = 16'd10;
        random_gaussian_normal[11] = 16'd341;
        random_gaussian_normal[12] = 16'd379;
        random_gaussian_normal[13] = 16'd138;
        random_gaussian_normal[14] = 16'd299;
        random_gaussian_normal[15] = 16'd401;
        random_gaussian_normal[16] = 16'd107;
        random_gaussian_normal[17] = 16'd442;
        random_gaussian_normal[18] = 16'd13;
        random_gaussian_normal[19] = 16'd55;
        random_gaussian_normal[20] = 16'd243;
        random_gaussian_normal[21] = 16'd46;
        random_gaussian_normal[22] = 16'd85;
        random_gaussian_normal[23] = 16'd153;
        random_gaussian_normal[24] = 16'd365;
        random_gaussian_normal[25] = 16'd72;
        random_gaussian_normal[26] = 16'd9;
        random_gaussian_normal[27] = 16'd109;
        random_gaussian_normal[28] = 16'd70;
        random_gaussian_normal[29] = 16'd217;
        random_gaussian_normal[30] = 16'd353;
        random_gaussian_normal[31] = 16'd87;
        random_gaussian_normal[32] = 16'd65;
        random_gaussian_normal[33] = 16'd286;
        random_gaussian_normal[34] = 16'd202;
        random_gaussian_normal[35] = 16'd244;
        random_gaussian_normal[36] = 16'd172;
        random_gaussian_normal[37] = 16'd120;
        random_gaussian_normal[38] = 16'd80;
        random_gaussian_normal[39] = 16'd91;
        random_gaussian_normal[40] = 16'd262;
        random_gaussian_normal[41] = 16'd499;
        random_gaussian_normal[42] = 16'd55;
        random_gaussian_normal[43] = 16'd133;
        random_gaussian_normal[44] = 16'd76;
        random_gaussian_normal[45] = 16'd45;
        random_gaussian_normal[46] = 16'd100;
        random_gaussian_normal[47] = 16'd172;
        random_gaussian_normal[48] = 16'd565;
        random_gaussian_normal[49] = 16'd217;
        random_gaussian_normal[50] = 16'd235;
        random_gaussian_normal[51] = 16'd4;
        random_gaussian_normal[52] = 16'd51;
        random_gaussian_normal[53] = 16'd34;
        random_gaussian_normal[54] = 16'd154;
        random_gaussian_normal[55] = 16'd369;
        random_gaussian_normal[56] = 16'd63;
        random_gaussian_normal[57] = 16'd57;
        random_gaussian_normal[58] = 16'd162;
        random_gaussian_normal[59] = 16'd400;
        random_gaussian_normal[60] = 16'd116;
        random_gaussian_normal[61] = 16'd85;
        random_gaussian_normal[62] = 16'd118;
        random_gaussian_normal[63] = 16'd216;
        random_gaussian_normal[64] = 16'd446;
        random_gaussian_normal[65] = 16'd254;
        random_gaussian_normal[66] = 16'd53;
        random_gaussian_normal[67] = 16'd404;
        random_gaussian_normal[68] = 16'd282;
        random_gaussian_normal[69] = 16'd183;
        random_gaussian_normal[70] = 16'd396;
        random_gaussian_normal[71] = 16'd124;
        random_gaussian_normal[72] = 16'd329;
        random_gaussian_normal[73] = 16'd109;
        random_gaussian_normal[74] = 16'd128;
        random_gaussian_normal[75] = 16'd176;
        random_gaussian_normal[76] = 16'd16;
        random_gaussian_normal[77] = 16'd131;
        random_gaussian_normal[78] = 16'd431;
        random_gaussian_normal[79] = 16'd102;
        random_gaussian_normal[80] = 16'd260;
        random_gaussian_normal[81] = 16'd411;
        random_gaussian_normal[82] = 16'd165;
        random_gaussian_normal[83] = 16'd95;
        random_gaussian_normal[84] = 16'd5;
        random_gaussian_normal[85] = 16'd159;
        random_gaussian_normal[86] = 16'd430;
        random_gaussian_normal[87] = 16'd223;
        random_gaussian_normal[88] = 16'd319;
        random_gaussian_normal[89] = 16'd608;
        random_gaussian_normal[90] = 16'd235;
        random_gaussian_normal[91] = 16'd58;
        random_gaussian_normal[92] = 16'd313;
        random_gaussian_normal[93] = 16'd64;
        random_gaussian_normal[94] = 16'd376;
        random_gaussian_normal[95] = 16'd19;
        random_gaussian_normal[96] = 16'd26;
        random_gaussian_normal[97] = 16'd374;
        random_gaussian_normal[98] = 16'd243;
        random_gaussian_normal[99] = 16'd182;
        random_gaussian_normal[100] = 16'd319;
        random_gaussian_normal[101] = 16'd325;
        random_gaussian_normal[102] = 16'd90;
        random_gaussian_normal[103] = 16'd68;
        random_gaussian_normal[104] = 16'd394;
        random_gaussian_normal[105] = 16'd40;
        random_gaussian_normal[106] = 16'd97;
        random_gaussian_normal[107] = 16'd278;
        random_gaussian_normal[108] = 16'd119;
        random_gaussian_normal[109] = 16'd292;
        random_gaussian_normal[110] = 16'd391;
        random_gaussian_normal[111] = 16'd526;
        random_gaussian_normal[112] = 16'd138;
        random_gaussian_normal[113] = 16'd95;
        random_gaussian_normal[114] = 16'd206;
        random_gaussian_normal[115] = 16'd120;
        random_gaussian_normal[116] = 16'd42;
        random_gaussian_normal[117] = 16'd403;
        random_gaussian_normal[118] = 16'd78;
        random_gaussian_normal[119] = 16'd347;
        random_gaussian_normal[120] = 16'd210;
        random_gaussian_normal[121] = 16'd239;
        random_gaussian_normal[122] = 16'd131;
        random_gaussian_normal[123] = 16'd149;
        random_gaussian_normal[124] = 16'd370;
        random_gaussian_normal[125] = 16'd321;
        random_gaussian_normal[126] = 16'd328;
        random_gaussian_normal[127] = 16'd267;
        random_gaussian_normal[128] = 16'd27;
        random_gaussian_normal[129] = 16'd1;
        random_gaussian_normal[130] = 16'd33;
        random_gaussian_normal[131] = 16'd410;
        random_gaussian_normal[132] = 16'd198;
        random_gaussian_normal[133] = 16'd5;
        random_gaussian_normal[134] = 16'd81;
        random_gaussian_normal[135] = 16'd284;
        random_gaussian_normal[136] = 16'd570;
        random_gaussian_normal[137] = 16'd26;
        random_gaussian_normal[138] = 16'd177;
        random_gaussian_normal[139] = 16'd284;
        random_gaussian_normal[140] = 16'd66;
        random_gaussian_normal[141] = 16'd154;
        random_gaussian_normal[142] = 16'd211;
        random_gaussian_normal[143] = 16'd240;
        random_gaussian_normal[144] = 16'd383;
        random_gaussian_normal[145] = 16'd555;
        random_gaussian_normal[146] = 16'd226;
        random_gaussian_normal[147] = 16'd237;
        random_gaussian_normal[148] = 16'd61;
        random_gaussian_normal[149] = 16'd80;
        random_gaussian_normal[150] = 16'd288;
        random_gaussian_normal[151] = 16'd389;
        random_gaussian_normal[152] = 16'd255;
        random_gaussian_normal[153] = 16'd293;
        random_gaussian_normal[154] = 16'd233;
        random_gaussian_normal[155] = 16'd53;
        random_gaussian_normal[156] = 16'd382;
        random_gaussian_normal[157] = 16'd28;
        random_gaussian_normal[158] = 16'd193;
        random_gaussian_normal[159] = 16'd223;
        random_gaussian_normal[160] = 16'd267;
        random_gaussian_normal[161] = 16'd196;
        random_gaussian_normal[162] = 16'd142;
        random_gaussian_normal[163] = 16'd153;
        random_gaussian_normal[164] = 16'd94;
        random_gaussian_normal[165] = 16'd69;
        random_gaussian_normal[166] = 16'd123;
        random_gaussian_normal[167] = 16'd279;
        random_gaussian_normal[168] = 16'd130;
        random_gaussian_normal[169] = 16'd153;
        random_gaussian_normal[170] = 16'd149;
        random_gaussian_normal[171] = 16'd64;
        random_gaussian_normal[172] = 16'd152;
        random_gaussian_normal[173] = 16'd64;
        random_gaussian_normal[174] = 16'd561;
        random_gaussian_normal[175] = 16'd129;
        random_gaussian_normal[176] = 16'd25;
        random_gaussian_normal[177] = 16'd534;
        random_gaussian_normal[178] = 16'd554;
        random_gaussian_normal[179] = 16'd124;
        random_gaussian_normal[180] = 16'd10;
        random_gaussian_normal[181] = 16'd65;
        random_gaussian_normal[182] = 16'd274;
        random_gaussian_normal[183] = 16'd276;
        random_gaussian_normal[184] = 16'd137;
        random_gaussian_normal[185] = 16'd233;
        random_gaussian_normal[186] = 16'd370;
        random_gaussian_normal[187] = 16'd298;
        random_gaussian_normal[188] = 16'd439;
        random_gaussian_normal[189] = 16'd538;
        random_gaussian_normal[190] = 16'd337;
        random_gaussian_normal[191] = 16'd206;
        random_gaussian_normal[192] = 16'd248;
        random_gaussian_normal[193] = 16'd566;
        random_gaussian_normal[194] = 16'd169;
        random_gaussian_normal[195] = 16'd84;
        random_gaussian_normal[196] = 16'd64;
        random_gaussian_normal[197] = 16'd537;
        random_gaussian_normal[198] = 16'd226;
        random_gaussian_normal[199] = 16'd95;
        random_gaussian_normal[200] = 16'd241;
        random_gaussian_normal[201] = 16'd642;
        random_gaussian_normal[202] = 16'd186;
        random_gaussian_normal[203] = 16'd214;
        random_gaussian_normal[204] = 16'd317;
        random_gaussian_normal[205] = 16'd62;
        random_gaussian_normal[206] = 16'd155;
        random_gaussian_normal[207] = 16'd512;
        random_gaussian_normal[208] = 16'd99;
        random_gaussian_normal[209] = 16'd9;
        random_gaussian_normal[210] = 16'd111;
        random_gaussian_normal[211] = 16'd302;
        random_gaussian_normal[212] = 16'd224;
        random_gaussian_normal[213] = 16'd32;
        random_gaussian_normal[214] = 16'd180;
        random_gaussian_normal[215] = 16'd234;
        random_gaussian_normal[216] = 16'd85;
        random_gaussian_normal[217] = 16'd30;
        random_gaussian_normal[218] = 16'd76;
        random_gaussian_normal[219] = 16'd780;
        random_gaussian_normal[220] = 16'd132;
        random_gaussian_normal[221] = 16'd137;
        random_gaussian_normal[222] = 16'd86;
        random_gaussian_normal[223] = 16'd504;
        random_gaussian_normal[224] = 16'd168;
        random_gaussian_normal[225] = 16'd15;
        random_gaussian_normal[226] = 16'd126;
        random_gaussian_normal[227] = 16'd59;
        random_gaussian_normal[228] = 16'd222;
        random_gaussian_normal[229] = 16'd73;
        random_gaussian_normal[230] = 16'd391;
        random_gaussian_normal[231] = 16'd3;
        random_gaussian_normal[232] = 16'd87;
        random_gaussian_normal[233] = 16'd319;
        random_gaussian_normal[234] = 16'd39;
        random_gaussian_normal[235] = 16'd70;
        random_gaussian_normal[236] = 16'd63;
        random_gaussian_normal[237] = 16'd396;
        random_gaussian_normal[238] = 16'd278;
        random_gaussian_normal[239] = 16'd257;
        random_gaussian_normal[240] = 16'd262;
        random_gaussian_normal[241] = 16'd494;
        random_gaussian_normal[242] = 16'd146;
        random_gaussian_normal[243] = 16'd66;
        random_gaussian_normal[244] = 16'd182;
        random_gaussian_normal[245] = 16'd23;
        random_gaussian_normal[246] = 16'd16;
        random_gaussian_normal[247] = 16'd365;
        random_gaussian_normal[248] = 16'd113;
        random_gaussian_normal[249] = 16'd56;
        random_gaussian_normal[250] = 16'd153;
        random_gaussian_normal[251] = 16'd314;
        random_gaussian_normal[252] = 16'd290;
        random_gaussian_normal[253] = 16'd150;
        random_gaussian_normal[254] = 16'd84;
        random_gaussian_normal[255] = 16'd416;
        random_gaussian_normal[256] = 16'd119;
        random_gaussian_normal[257] = 16'd23;
        random_gaussian_normal[258] = 16'd623;
        random_gaussian_normal[259] = 16'd372;
        random_gaussian_normal[260] = 16'd192;
        random_gaussian_normal[261] = 16'd268;
        random_gaussian_normal[262] = 16'd97;
        random_gaussian_normal[263] = 16'd122;
        random_gaussian_normal[264] = 16'd318;
        random_gaussian_normal[265] = 16'd359;
        random_gaussian_normal[266] = 16'd182;
        random_gaussian_normal[267] = 16'd69;
        random_gaussian_normal[268] = 16'd204;
        random_gaussian_normal[269] = 16'd182;
        random_gaussian_normal[270] = 16'd234;
        random_gaussian_normal[271] = 16'd91;
        random_gaussian_normal[272] = 16'd9;
        random_gaussian_normal[273] = 16'd579;
        random_gaussian_normal[274] = 16'd319;
        random_gaussian_normal[275] = 16'd228;
        random_gaussian_normal[276] = 16'd82;
        random_gaussian_normal[277] = 16'd344;
        random_gaussian_normal[278] = 16'd279;
        random_gaussian_normal[279] = 16'd278;
        random_gaussian_normal[280] = 16'd118;
        random_gaussian_normal[281] = 16'd263;
        random_gaussian_normal[282] = 16'd439;
        random_gaussian_normal[283] = 16'd46;
        random_gaussian_normal[284] = 16'd184;
        random_gaussian_normal[285] = 16'd111;
        random_gaussian_normal[286] = 16'd189;
        random_gaussian_normal[287] = 16'd392;
        random_gaussian_normal[288] = 16'd328;
        random_gaussian_normal[289] = 16'd118;
        random_gaussian_normal[290] = 16'd86;
        random_gaussian_normal[291] = 16'd39;
        random_gaussian_normal[292] = 16'd108;
        random_gaussian_normal[293] = 16'd3;
        random_gaussian_normal[294] = 16'd274;
        random_gaussian_normal[295] = 16'd566;
        random_gaussian_normal[296] = 16'd299;
        random_gaussian_normal[297] = 16'd343;
        random_gaussian_normal[298] = 16'd321;
        random_gaussian_normal[299] = 16'd282;
        random_gaussian_normal[300] = 16'd90;
        random_gaussian_normal[301] = 16'd361;
        random_gaussian_normal[302] = 16'd619;
        random_gaussian_normal[303] = 16'd377;
        random_gaussian_normal[304] = 16'd4;
        random_gaussian_normal[305] = 16'd92;
        random_gaussian_normal[306] = 16'd112;
        random_gaussian_normal[307] = 16'd266;
        random_gaussian_normal[308] = 16'd263;
        random_gaussian_normal[309] = 16'd60;
        random_gaussian_normal[310] = 16'd241;
        random_gaussian_normal[311] = 16'd322;
        random_gaussian_normal[312] = 16'd133;
        random_gaussian_normal[313] = 16'd632;
        random_gaussian_normal[314] = 16'd55;
        random_gaussian_normal[315] = 16'd435;
        random_gaussian_normal[316] = 16'd483;
        random_gaussian_normal[317] = 16'd130;
        random_gaussian_normal[318] = 16'd127;
        random_gaussian_normal[319] = 16'd4;
        random_gaussian_normal[320] = 16'd465;
        random_gaussian_normal[321] = 16'd236;
        random_gaussian_normal[322] = 16'd126;
        random_gaussian_normal[323] = 16'd135;
        random_gaussian_normal[324] = 16'd17;
        random_gaussian_normal[325] = 16'd645;
        random_gaussian_normal[326] = 16'd42;
        random_gaussian_normal[327] = 16'd108;
        random_gaussian_normal[328] = 16'd114;
        random_gaussian_normal[329] = 16'd33;
        random_gaussian_normal[330] = 16'd162;
        random_gaussian_normal[331] = 16'd130;
        random_gaussian_normal[332] = 16'd30;
        random_gaussian_normal[333] = 16'd282;
        random_gaussian_normal[334] = 16'd145;
        random_gaussian_normal[335] = 16'd487;
        random_gaussian_normal[336] = 16'd457;
        random_gaussian_normal[337] = 16'd262;
        random_gaussian_normal[338] = 16'd289;
        random_gaussian_normal[339] = 16'd7;
        random_gaussian_normal[340] = 16'd162;
        random_gaussian_normal[341] = 16'd50;
        random_gaussian_normal[342] = 16'd42;
        random_gaussian_normal[343] = 16'd163;
        random_gaussian_normal[344] = 16'd59;
        random_gaussian_normal[345] = 16'd10;
        random_gaussian_normal[346] = 16'd13;
        random_gaussian_normal[347] = 16'd257;
        random_gaussian_normal[348] = 16'd92;
        random_gaussian_normal[349] = 16'd141;
        random_gaussian_normal[350] = 16'd347;
        random_gaussian_normal[351] = 16'd439;
        random_gaussian_normal[352] = 16'd65;
        random_gaussian_normal[353] = 16'd91;
        random_gaussian_normal[354] = 16'd312;
        random_gaussian_normal[355] = 16'd119;
        random_gaussian_normal[356] = 16'd40;
        random_gaussian_normal[357] = 16'd264;
        random_gaussian_normal[358] = 16'd74;
        random_gaussian_normal[359] = 16'd238;
        random_gaussian_normal[360] = 16'd34;
        random_gaussian_normal[361] = 16'd508;
        random_gaussian_normal[362] = 16'd233;
        random_gaussian_normal[363] = 16'd58;
        random_gaussian_normal[364] = 16'd214;
        random_gaussian_normal[365] = 16'd9;
        random_gaussian_normal[366] = 16'd201;
        random_gaussian_normal[367] = 16'd249;
        random_gaussian_normal[368] = 16'd255;
        random_gaussian_normal[369] = 16'd222;
        random_gaussian_normal[370] = 16'd140;
        random_gaussian_normal[371] = 16'd173;
        random_gaussian_normal[372] = 16'd150;
        random_gaussian_normal[373] = 16'd254;
        random_gaussian_normal[374] = 16'd269;
        random_gaussian_normal[375] = 16'd170;
        random_gaussian_normal[376] = 16'd259;
        random_gaussian_normal[377] = 16'd300;
        random_gaussian_normal[378] = 16'd189;
        random_gaussian_normal[379] = 16'd166;
        random_gaussian_normal[380] = 16'd307;
        random_gaussian_normal[381] = 16'd570;
        random_gaussian_normal[382] = 16'd207;
        random_gaussian_normal[383] = 16'd216;
        random_gaussian_normal[384] = 16'd178;
        random_gaussian_normal[385] = 16'd216;
        random_gaussian_normal[386] = 16'd289;
        random_gaussian_normal[387] = 16'd91;
        random_gaussian_normal[388] = 16'd271;
        random_gaussian_normal[389] = 16'd144;
        random_gaussian_normal[390] = 16'd376;
        random_gaussian_normal[391] = 16'd132;
        random_gaussian_normal[392] = 16'd379;
        random_gaussian_normal[393] = 16'd47;
        random_gaussian_normal[394] = 16'd82;
        random_gaussian_normal[395] = 16'd156;
        random_gaussian_normal[396] = 16'd37;
        random_gaussian_normal[397] = 16'd227;
        random_gaussian_normal[398] = 16'd124;
        random_gaussian_normal[399] = 16'd138;
        random_gaussian_normal[400] = 16'd406;
        random_gaussian_normal[401] = 16'd24;
        random_gaussian_normal[402] = 16'd139;
        random_gaussian_normal[403] = 16'd31;
        random_gaussian_normal[404] = 16'd92;
        random_gaussian_normal[405] = 16'd164;
        random_gaussian_normal[406] = 16'd152;
        random_gaussian_normal[407] = 16'd30;
        random_gaussian_normal[408] = 16'd212;
        random_gaussian_normal[409] = 16'd92;
        random_gaussian_normal[410] = 16'd99;
        random_gaussian_normal[411] = 16'd281;
        random_gaussian_normal[412] = 16'd7;
        random_gaussian_normal[413] = 16'd331;
        random_gaussian_normal[414] = 16'd405;
        random_gaussian_normal[415] = 16'd765;
        random_gaussian_normal[416] = 16'd63;
        random_gaussian_normal[417] = 16'd105;
        random_gaussian_normal[418] = 16'd212;
        random_gaussian_normal[419] = 16'd53;
        random_gaussian_normal[420] = 16'd274;
        random_gaussian_normal[421] = 16'd184;
        random_gaussian_normal[422] = 16'd245;
        random_gaussian_normal[423] = 16'd85;
        random_gaussian_normal[424] = 16'd133;
        random_gaussian_normal[425] = 16'd255;
        random_gaussian_normal[426] = 16'd106;
        random_gaussian_normal[427] = 16'd48;
        random_gaussian_normal[428] = 16'd227;
        random_gaussian_normal[429] = 16'd196;
        random_gaussian_normal[430] = 16'd184;
        random_gaussian_normal[431] = 16'd374;
        random_gaussian_normal[432] = 16'd55;
        random_gaussian_normal[433] = 16'd487;
        random_gaussian_normal[434] = 16'd401;
        random_gaussian_normal[435] = 16'd533;
        random_gaussian_normal[436] = 16'd367;
        random_gaussian_normal[437] = 16'd502;
        random_gaussian_normal[438] = 16'd31;
        random_gaussian_normal[439] = 16'd324;
        random_gaussian_normal[440] = 16'd110;
        random_gaussian_normal[441] = 16'd81;
        random_gaussian_normal[442] = 16'd56;
        random_gaussian_normal[443] = 16'd49;
        random_gaussian_normal[444] = 16'd348;
        random_gaussian_normal[445] = 16'd46;
        random_gaussian_normal[446] = 16'd266;
        random_gaussian_normal[447] = 16'd185;
        random_gaussian_normal[448] = 16'd481;
        random_gaussian_normal[449] = 16'd34;
        random_gaussian_normal[450] = 16'd164;
        random_gaussian_normal[451] = 16'd422;
        random_gaussian_normal[452] = 16'd63;
        random_gaussian_normal[453] = 16'd178;
        random_gaussian_normal[454] = 16'd681;
        random_gaussian_normal[455] = 16'd161;
        random_gaussian_normal[456] = 16'd333;
        random_gaussian_normal[457] = 16'd165;
        random_gaussian_normal[458] = 16'd224;
        random_gaussian_normal[459] = 16'd325;
        random_gaussian_normal[460] = 16'd151;
        random_gaussian_normal[461] = 16'd385;
        random_gaussian_normal[462] = 16'd58;
        random_gaussian_normal[463] = 16'd400;
        random_gaussian_normal[464] = 16'd518;
        random_gaussian_normal[465] = 16'd47;
        random_gaussian_normal[466] = 16'd155;
        random_gaussian_normal[467] = 16'd180;
        random_gaussian_normal[468] = 16'd421;
        random_gaussian_normal[469] = 16'd35;
        random_gaussian_normal[470] = 16'd129;
        random_gaussian_normal[471] = 16'd400;
        random_gaussian_normal[472] = 16'd114;
        random_gaussian_normal[473] = 16'd551;
        random_gaussian_normal[474] = 16'd247;
        random_gaussian_normal[475] = 16'd94;
        random_gaussian_normal[476] = 16'd162;
        random_gaussian_normal[477] = 16'd103;
        random_gaussian_normal[478] = 16'd152;
        random_gaussian_normal[479] = 16'd328;
        random_gaussian_normal[480] = 16'd16;
        random_gaussian_normal[481] = 16'd274;
        random_gaussian_normal[482] = 16'd4;
        random_gaussian_normal[483] = 16'd14;
        random_gaussian_normal[484] = 16'd8;
        random_gaussian_normal[485] = 16'd121;
        random_gaussian_normal[486] = 16'd317;
        random_gaussian_normal[487] = 16'd437;
        random_gaussian_normal[488] = 16'd202;
        random_gaussian_normal[489] = 16'd16;
        random_gaussian_normal[490] = 16'd191;
        random_gaussian_normal[491] = 16'd14;
        random_gaussian_normal[492] = 16'd103;
        random_gaussian_normal[493] = 16'd242;
        random_gaussian_normal[494] = 16'd136;
        random_gaussian_normal[495] = 16'd105;
        random_gaussian_normal[496] = 16'd268;
        random_gaussian_normal[497] = 16'd115;
        random_gaussian_normal[498] = 16'd472;
        random_gaussian_normal[499] = 16'd15;
        random_gaussian_normal[500] = 16'd104;
        random_gaussian_normal[501] = 16'd356;
        random_gaussian_normal[502] = 16'd75;
        random_gaussian_normal[503] = 16'd16;
        random_gaussian_normal[504] = 16'd225;
        random_gaussian_normal[505] = 16'd359;
        random_gaussian_normal[506] = 16'd666;
        random_gaussian_normal[507] = 16'd159;
        random_gaussian_normal[508] = 16'd67;
        random_gaussian_normal[509] = 16'd109;
        random_gaussian_normal[510] = 16'd242;
        random_gaussian_normal[511] = 16'd327;
        random_gaussian_normal[512] = 16'd137;
        random_gaussian_normal[513] = 16'd410;
        random_gaussian_normal[514] = 16'd240;
        random_gaussian_normal[515] = 16'd145;
        random_gaussian_normal[516] = 16'd131;
        random_gaussian_normal[517] = 16'd494;
        random_gaussian_normal[518] = 16'd270;
        random_gaussian_normal[519] = 16'd191;
        random_gaussian_normal[520] = 16'd181;
        random_gaussian_normal[521] = 16'd495;
        random_gaussian_normal[522] = 16'd59;
        random_gaussian_normal[523] = 16'd43;
        random_gaussian_normal[524] = 16'd188;
        random_gaussian_normal[525] = 16'd210;
        random_gaussian_normal[526] = 16'd82;
        random_gaussian_normal[527] = 16'd144;
        random_gaussian_normal[528] = 16'd88;
        random_gaussian_normal[529] = 16'd87;
        random_gaussian_normal[530] = 16'd276;
        random_gaussian_normal[531] = 16'd276;
        random_gaussian_normal[532] = 16'd84;
        random_gaussian_normal[533] = 16'd250;
        random_gaussian_normal[534] = 16'd336;
        random_gaussian_normal[535] = 16'd88;
        random_gaussian_normal[536] = 16'd23;
        random_gaussian_normal[537] = 16'd65;
        random_gaussian_normal[538] = 16'd99;
        random_gaussian_normal[539] = 16'd48;
        random_gaussian_normal[540] = 16'd559;
        random_gaussian_normal[541] = 16'd91;
        random_gaussian_normal[542] = 16'd158;
        random_gaussian_normal[543] = 16'd13;
        random_gaussian_normal[544] = 16'd348;
        random_gaussian_normal[545] = 16'd210;
        random_gaussian_normal[546] = 16'd188;
        random_gaussian_normal[547] = 16'd2;
        random_gaussian_normal[548] = 16'd176;
        random_gaussian_normal[549] = 16'd317;
        random_gaussian_normal[550] = 16'd476;
        random_gaussian_normal[551] = 16'd274;
        random_gaussian_normal[552] = 16'd133;
        random_gaussian_normal[553] = 16'd379;
        random_gaussian_normal[554] = 16'd302;
        random_gaussian_normal[555] = 16'd491;
        random_gaussian_normal[556] = 16'd165;
        random_gaussian_normal[557] = 16'd388;
        random_gaussian_normal[558] = 16'd156;
        random_gaussian_normal[559] = 16'd486;
        random_gaussian_normal[560] = 16'd91;
        random_gaussian_normal[561] = 16'd71;
        random_gaussian_normal[562] = 16'd266;
        random_gaussian_normal[563] = 16'd295;
        random_gaussian_normal[564] = 16'd28;
        random_gaussian_normal[565] = 16'd291;
        random_gaussian_normal[566] = 16'd231;
        random_gaussian_normal[567] = 16'd257;
        random_gaussian_normal[568] = 16'd205;
        random_gaussian_normal[569] = 16'd421;
        random_gaussian_normal[570] = 16'd245;
        random_gaussian_normal[571] = 16'd152;
        random_gaussian_normal[572] = 16'd427;
        random_gaussian_normal[573] = 16'd218;
        random_gaussian_normal[574] = 16'd24;
        random_gaussian_normal[575] = 16'd129;
        random_gaussian_normal[576] = 16'd50;
        random_gaussian_normal[577] = 16'd25;
        random_gaussian_normal[578] = 16'd558;
        random_gaussian_normal[579] = 16'd294;
        random_gaussian_normal[580] = 16'd329;
        random_gaussian_normal[581] = 16'd107;
        random_gaussian_normal[582] = 16'd24;
        random_gaussian_normal[583] = 16'd68;
        random_gaussian_normal[584] = 16'd152;
        random_gaussian_normal[585] = 16'd11;
        random_gaussian_normal[586] = 16'd164;
        random_gaussian_normal[587] = 16'd260;
        random_gaussian_normal[588] = 16'd184;
        random_gaussian_normal[589] = 16'd149;
        random_gaussian_normal[590] = 16'd260;
        random_gaussian_normal[591] = 16'd443;
        random_gaussian_normal[592] = 16'd64;
        random_gaussian_normal[593] = 16'd534;
        random_gaussian_normal[594] = 16'd634;
        random_gaussian_normal[595] = 16'd216;
        random_gaussian_normal[596] = 16'd301;
        random_gaussian_normal[597] = 16'd485;
        random_gaussian_normal[598] = 16'd272;
        random_gaussian_normal[599] = 16'd83;
        random_gaussian_normal[600] = 16'd184;
        random_gaussian_normal[601] = 16'd39;
        random_gaussian_normal[602] = 16'd189;
        random_gaussian_normal[603] = 16'd790;
        random_gaussian_normal[604] = 16'd77;
        random_gaussian_normal[605] = 16'd138;
        random_gaussian_normal[606] = 16'd7;
        random_gaussian_normal[607] = 16'd41;
        random_gaussian_normal[608] = 16'd110;
        random_gaussian_normal[609] = 16'd164;
        random_gaussian_normal[610] = 16'd227;
        random_gaussian_normal[611] = 16'd18;
        random_gaussian_normal[612] = 16'd235;
        random_gaussian_normal[613] = 16'd352;
        random_gaussian_normal[614] = 16'd340;
        random_gaussian_normal[615] = 16'd179;
        random_gaussian_normal[616] = 16'd125;
        random_gaussian_normal[617] = 16'd67;
        random_gaussian_normal[618] = 16'd225;
        random_gaussian_normal[619] = 16'd166;
        random_gaussian_normal[620] = 16'd130;
        random_gaussian_normal[621] = 16'd217;
        random_gaussian_normal[622] = 16'd636;
        random_gaussian_normal[623] = 16'd78;
        random_gaussian_normal[624] = 16'd331;
        random_gaussian_normal[625] = 16'd160;
        random_gaussian_normal[626] = 16'd10;
        random_gaussian_normal[627] = 16'd112;
        random_gaussian_normal[628] = 16'd104;
        random_gaussian_normal[629] = 16'd601;
        random_gaussian_normal[630] = 16'd198;
        random_gaussian_normal[631] = 16'd1;
        random_gaussian_normal[632] = 16'd171;
        random_gaussian_normal[633] = 16'd545;
        random_gaussian_normal[634] = 16'd225;
        random_gaussian_normal[635] = 16'd188;
        random_gaussian_normal[636] = 16'd69;
        random_gaussian_normal[637] = 16'd568;
        random_gaussian_normal[638] = 16'd471;
        random_gaussian_normal[639] = 16'd325;
        random_gaussian_normal[640] = 16'd69;
        random_gaussian_normal[641] = 16'd73;
        random_gaussian_normal[642] = 16'd122;
        random_gaussian_normal[643] = 16'd20;
        random_gaussian_normal[644] = 16'd3;
        random_gaussian_normal[645] = 16'd237;
        random_gaussian_normal[646] = 16'd239;
        random_gaussian_normal[647] = 16'd370;
        random_gaussian_normal[648] = 16'd85;
        random_gaussian_normal[649] = 16'd25;
        random_gaussian_normal[650] = 16'd400;
        random_gaussian_normal[651] = 16'd65;
        random_gaussian_normal[652] = 16'd74;
        random_gaussian_normal[653] = 16'd304;
        random_gaussian_normal[654] = 16'd175;
        random_gaussian_normal[655] = 16'd395;
        random_gaussian_normal[656] = 16'd117;
        random_gaussian_normal[657] = 16'd198;
        random_gaussian_normal[658] = 16'd7;
        random_gaussian_normal[659] = 16'd354;
        random_gaussian_normal[660] = 16'd146;
        random_gaussian_normal[661] = 16'd272;
        random_gaussian_normal[662] = 16'd128;
        random_gaussian_normal[663] = 16'd162;
        random_gaussian_normal[664] = 16'd472;
        random_gaussian_normal[665] = 16'd40;
        random_gaussian_normal[666] = 16'd347;
        random_gaussian_normal[667] = 16'd211;
        random_gaussian_normal[668] = 16'd69;
        random_gaussian_normal[669] = 16'd166;
        random_gaussian_normal[670] = 16'd88;
        random_gaussian_normal[671] = 16'd60;
        random_gaussian_normal[672] = 16'd176;
        random_gaussian_normal[673] = 16'd60;
        random_gaussian_normal[674] = 16'd33;
        random_gaussian_normal[675] = 16'd247;
        random_gaussian_normal[676] = 16'd79;
        random_gaussian_normal[677] = 16'd153;
        random_gaussian_normal[678] = 16'd18;
        random_gaussian_normal[679] = 16'd84;
        random_gaussian_normal[680] = 16'd340;
        random_gaussian_normal[681] = 16'd273;
        random_gaussian_normal[682] = 16'd36;
        random_gaussian_normal[683] = 16'd127;
        random_gaussian_normal[684] = 16'd53;
        random_gaussian_normal[685] = 16'd26;
        random_gaussian_normal[686] = 16'd137;
        random_gaussian_normal[687] = 16'd108;
        random_gaussian_normal[688] = 16'd90;
        random_gaussian_normal[689] = 16'd98;
        random_gaussian_normal[690] = 16'd42;
        random_gaussian_normal[691] = 16'd30;
        random_gaussian_normal[692] = 16'd311;
        random_gaussian_normal[693] = 16'd342;
        random_gaussian_normal[694] = 16'd32;
        random_gaussian_normal[695] = 16'd544;
        random_gaussian_normal[696] = 16'd100;
        random_gaussian_normal[697] = 16'd402;
        random_gaussian_normal[698] = 16'd85;
        random_gaussian_normal[699] = 16'd157;
        random_gaussian_normal[700] = 16'd98;
        random_gaussian_normal[701] = 16'd302;
        random_gaussian_normal[702] = 16'd7;
        random_gaussian_normal[703] = 16'd47;
        random_gaussian_normal[704] = 16'd27;
        random_gaussian_normal[705] = 16'd778;
        random_gaussian_normal[706] = 16'd185;
        random_gaussian_normal[707] = 16'd308;
        random_gaussian_normal[708] = 16'd15;
        random_gaussian_normal[709] = 16'd227;
        random_gaussian_normal[710] = 16'd137;
        random_gaussian_normal[711] = 16'd247;
        random_gaussian_normal[712] = 16'd34;
        random_gaussian_normal[713] = 16'd265;
        random_gaussian_normal[714] = 16'd175;
        random_gaussian_normal[715] = 16'd467;
        random_gaussian_normal[716] = 16'd233;
        random_gaussian_normal[717] = 16'd374;
        random_gaussian_normal[718] = 16'd203;
        random_gaussian_normal[719] = 16'd67;
        random_gaussian_normal[720] = 16'd172;
        random_gaussian_normal[721] = 16'd23;
        random_gaussian_normal[722] = 16'd400;
        random_gaussian_normal[723] = 16'd243;
        random_gaussian_normal[724] = 16'd253;
        random_gaussian_normal[725] = 16'd87;
        random_gaussian_normal[726] = 16'd403;
        random_gaussian_normal[727] = 16'd100;
        random_gaussian_normal[728] = 16'd308;
        random_gaussian_normal[729] = 16'd182;
        random_gaussian_normal[730] = 16'd513;
        random_gaussian_normal[731] = 16'd311;
        random_gaussian_normal[732] = 16'd6;
        random_gaussian_normal[733] = 16'd62;
        random_gaussian_normal[734] = 16'd20;
        random_gaussian_normal[735] = 16'd393;
        random_gaussian_normal[736] = 16'd257;
        random_gaussian_normal[737] = 16'd26;
        random_gaussian_normal[738] = 16'd122;
        random_gaussian_normal[739] = 16'd128;
        random_gaussian_normal[740] = 16'd351;
        random_gaussian_normal[741] = 16'd448;
        random_gaussian_normal[742] = 16'd408;
        random_gaussian_normal[743] = 16'd3;
        random_gaussian_normal[744] = 16'd502;
        random_gaussian_normal[745] = 16'd255;
        random_gaussian_normal[746] = 16'd37;
        random_gaussian_normal[747] = 16'd294;
        random_gaussian_normal[748] = 16'd123;
        random_gaussian_normal[749] = 16'd7;
        random_gaussian_normal[750] = 16'd122;
        random_gaussian_normal[751] = 16'd182;
        random_gaussian_normal[752] = 16'd26;
        random_gaussian_normal[753] = 16'd452;
        random_gaussian_normal[754] = 16'd6;
        random_gaussian_normal[755] = 16'd430;
        random_gaussian_normal[756] = 16'd280;
        random_gaussian_normal[757] = 16'd36;
        random_gaussian_normal[758] = 16'd119;
        random_gaussian_normal[759] = 16'd450;
        random_gaussian_normal[760] = 16'd239;
        random_gaussian_normal[761] = 16'd90;
        random_gaussian_normal[762] = 16'd128;
        random_gaussian_normal[763] = 16'd171;
        random_gaussian_normal[764] = 16'd167;
        random_gaussian_normal[765] = 16'd4;
        random_gaussian_normal[766] = 16'd444;
        random_gaussian_normal[767] = 16'd15;
        random_gaussian_normal[768] = 16'd532;
        random_gaussian_normal[769] = 16'd314;
        random_gaussian_normal[770] = 16'd129;
        random_gaussian_normal[771] = 16'd235;
        random_gaussian_normal[772] = 16'd130;
        random_gaussian_normal[773] = 16'd23;
        random_gaussian_normal[774] = 16'd115;
        random_gaussian_normal[775] = 16'd808;
        random_gaussian_normal[776] = 16'd0;
        random_gaussian_normal[777] = 16'd30;
        random_gaussian_normal[778] = 16'd485;
        random_gaussian_normal[779] = 16'd154;
        random_gaussian_normal[780] = 16'd5;
        random_gaussian_normal[781] = 16'd97;
        random_gaussian_normal[782] = 16'd338;
        random_gaussian_normal[783] = 16'd56;
        random_gaussian_normal[784] = 16'd71;
        random_gaussian_normal[785] = 16'd53;
        random_gaussian_normal[786] = 16'd47;
        random_gaussian_normal[787] = 16'd79;
        random_gaussian_normal[788] = 16'd127;
        random_gaussian_normal[789] = 16'd381;
        random_gaussian_normal[790] = 16'd263;
        random_gaussian_normal[791] = 16'd297;
        random_gaussian_normal[792] = 16'd254;
        random_gaussian_normal[793] = 16'd0;
        random_gaussian_normal[794] = 16'd270;
        random_gaussian_normal[795] = 16'd277;
        random_gaussian_normal[796] = 16'd176;
        random_gaussian_normal[797] = 16'd222;
        random_gaussian_normal[798] = 16'd313;
        random_gaussian_normal[799] = 16'd305;
        random_gaussian_normal[800] = 16'd373;
        random_gaussian_normal[801] = 16'd105;
        random_gaussian_normal[802] = 16'd141;
        random_gaussian_normal[803] = 16'd144;
        random_gaussian_normal[804] = 16'd229;
        random_gaussian_normal[805] = 16'd104;
        random_gaussian_normal[806] = 16'd258;
        random_gaussian_normal[807] = 16'd338;
        random_gaussian_normal[808] = 16'd142;
        random_gaussian_normal[809] = 16'd219;
        random_gaussian_normal[810] = 16'd32;
        random_gaussian_normal[811] = 16'd62;
        random_gaussian_normal[812] = 16'd44;
        random_gaussian_normal[813] = 16'd9;
        random_gaussian_normal[814] = 16'd163;
        random_gaussian_normal[815] = 16'd253;
        random_gaussian_normal[816] = 16'd107;
        random_gaussian_normal[817] = 16'd214;
        random_gaussian_normal[818] = 16'd60;
        random_gaussian_normal[819] = 16'd393;
        random_gaussian_normal[820] = 16'd33;
        random_gaussian_normal[821] = 16'd15;
        random_gaussian_normal[822] = 16'd504;
        random_gaussian_normal[823] = 16'd190;
        random_gaussian_normal[824] = 16'd185;
        random_gaussian_normal[825] = 16'd151;
        random_gaussian_normal[826] = 16'd337;
        random_gaussian_normal[827] = 16'd421;
        random_gaussian_normal[828] = 16'd88;
        random_gaussian_normal[829] = 16'd107;
        random_gaussian_normal[830] = 16'd357;
        random_gaussian_normal[831] = 16'd46;
        random_gaussian_normal[832] = 16'd414;
        random_gaussian_normal[833] = 16'd81;
        random_gaussian_normal[834] = 16'd62;
        random_gaussian_normal[835] = 16'd118;
        random_gaussian_normal[836] = 16'd76;
        random_gaussian_normal[837] = 16'd173;
        random_gaussian_normal[838] = 16'd123;
        random_gaussian_normal[839] = 16'd532;
        random_gaussian_normal[840] = 16'd311;
        random_gaussian_normal[841] = 16'd106;
        random_gaussian_normal[842] = 16'd128;
        random_gaussian_normal[843] = 16'd56;
        random_gaussian_normal[844] = 16'd73;
        random_gaussian_normal[845] = 16'd194;
        random_gaussian_normal[846] = 16'd64;
        random_gaussian_normal[847] = 16'd163;
        random_gaussian_normal[848] = 16'd146;
        random_gaussian_normal[849] = 16'd211;
        random_gaussian_normal[850] = 16'd341;
        random_gaussian_normal[851] = 16'd68;
        random_gaussian_normal[852] = 16'd45;
        random_gaussian_normal[853] = 16'd226;
        random_gaussian_normal[854] = 16'd303;
        random_gaussian_normal[855] = 16'd163;
        random_gaussian_normal[856] = 16'd33;
        random_gaussian_normal[857] = 16'd82;
        random_gaussian_normal[858] = 16'd67;
        random_gaussian_normal[859] = 16'd300;
        random_gaussian_normal[860] = 16'd90;
        random_gaussian_normal[861] = 16'd86;
        random_gaussian_normal[862] = 16'd39;
        random_gaussian_normal[863] = 16'd474;
        random_gaussian_normal[864] = 16'd125;
        random_gaussian_normal[865] = 16'd249;
        random_gaussian_normal[866] = 16'd501;
        random_gaussian_normal[867] = 16'd4;
        random_gaussian_normal[868] = 16'd464;
        random_gaussian_normal[869] = 16'd152;
        random_gaussian_normal[870] = 16'd217;
        random_gaussian_normal[871] = 16'd115;
        random_gaussian_normal[872] = 16'd16;
        random_gaussian_normal[873] = 16'd141;
        random_gaussian_normal[874] = 16'd283;
        random_gaussian_normal[875] = 16'd97;
        random_gaussian_normal[876] = 16'd465;
        random_gaussian_normal[877] = 16'd474;
        random_gaussian_normal[878] = 16'd205;
        random_gaussian_normal[879] = 16'd280;
        random_gaussian_normal[880] = 16'd690;
        random_gaussian_normal[881] = 16'd253;
        random_gaussian_normal[882] = 16'd576;
        random_gaussian_normal[883] = 16'd121;
        random_gaussian_normal[884] = 16'd36;
        random_gaussian_normal[885] = 16'd119;
        random_gaussian_normal[886] = 16'd56;
        random_gaussian_normal[887] = 16'd65;
        random_gaussian_normal[888] = 16'd91;
        random_gaussian_normal[889] = 16'd239;
        random_gaussian_normal[890] = 16'd287;
        random_gaussian_normal[891] = 16'd79;
        random_gaussian_normal[892] = 16'd86;
        random_gaussian_normal[893] = 16'd39;
        random_gaussian_normal[894] = 16'd8;
        random_gaussian_normal[895] = 16'd182;
        random_gaussian_normal[896] = 16'd111;
        random_gaussian_normal[897] = 16'd233;
        random_gaussian_normal[898] = 16'd96;
        random_gaussian_normal[899] = 16'd9;
        random_gaussian_normal[900] = 16'd4;
        random_gaussian_normal[901] = 16'd196;
        random_gaussian_normal[902] = 16'd93;
        random_gaussian_normal[903] = 16'd267;
        random_gaussian_normal[904] = 16'd173;
        random_gaussian_normal[905] = 16'd249;
        random_gaussian_normal[906] = 16'd188;
        random_gaussian_normal[907] = 16'd5;
        random_gaussian_normal[908] = 16'd94;
        random_gaussian_normal[909] = 16'd64;
        random_gaussian_normal[910] = 16'd203;
        random_gaussian_normal[911] = 16'd109;
        random_gaussian_normal[912] = 16'd292;
        random_gaussian_normal[913] = 16'd259;
        random_gaussian_normal[914] = 16'd99;
        random_gaussian_normal[915] = 16'd646;
        random_gaussian_normal[916] = 16'd256;
        random_gaussian_normal[917] = 16'd462;
        random_gaussian_normal[918] = 16'd127;
        random_gaussian_normal[919] = 16'd5;
        random_gaussian_normal[920] = 16'd198;
        random_gaussian_normal[921] = 16'd601;
        random_gaussian_normal[922] = 16'd117;
        random_gaussian_normal[923] = 16'd116;
        random_gaussian_normal[924] = 16'd135;
        random_gaussian_normal[925] = 16'd73;
        random_gaussian_normal[926] = 16'd522;
        random_gaussian_normal[927] = 16'd321;
        random_gaussian_normal[928] = 16'd442;
        random_gaussian_normal[929] = 16'd96;
        random_gaussian_normal[930] = 16'd287;
        random_gaussian_normal[931] = 16'd529;
        random_gaussian_normal[932] = 16'd385;
        random_gaussian_normal[933] = 16'd209;
        random_gaussian_normal[934] = 16'd178;
        random_gaussian_normal[935] = 16'd308;
        random_gaussian_normal[936] = 16'd167;
        random_gaussian_normal[937] = 16'd13;
        random_gaussian_normal[938] = 16'd71;
        random_gaussian_normal[939] = 16'd55;
        random_gaussian_normal[940] = 16'd449;
        random_gaussian_normal[941] = 16'd110;
        random_gaussian_normal[942] = 16'd181;
        random_gaussian_normal[943] = 16'd35;
        random_gaussian_normal[944] = 16'd291;
        random_gaussian_normal[945] = 16'd29;
        random_gaussian_normal[946] = 16'd66;
        random_gaussian_normal[947] = 16'd457;
        random_gaussian_normal[948] = 16'd459;
        random_gaussian_normal[949] = 16'd176;
        random_gaussian_normal[950] = 16'd100;
        random_gaussian_normal[951] = 16'd171;
        random_gaussian_normal[952] = 16'd95;
        random_gaussian_normal[953] = 16'd122;
        random_gaussian_normal[954] = 16'd90;
        random_gaussian_normal[955] = 16'd249;
        random_gaussian_normal[956] = 16'd52;
        random_gaussian_normal[957] = 16'd174;
        random_gaussian_normal[958] = 16'd173;
        random_gaussian_normal[959] = 16'd228;
        random_gaussian_normal[960] = 16'd146;
        random_gaussian_normal[961] = 16'd338;
        random_gaussian_normal[962] = 16'd412;
        random_gaussian_normal[963] = 16'd333;
        random_gaussian_normal[964] = 16'd503;
        random_gaussian_normal[965] = 16'd1;
        random_gaussian_normal[966] = 16'd85;
        random_gaussian_normal[967] = 16'd507;
        random_gaussian_normal[968] = 16'd183;
        random_gaussian_normal[969] = 16'd257;
        random_gaussian_normal[970] = 16'd145;
        random_gaussian_normal[971] = 16'd39;
        random_gaussian_normal[972] = 16'd451;
        random_gaussian_normal[973] = 16'd355;
        random_gaussian_normal[974] = 16'd35;
        random_gaussian_normal[975] = 16'd220;
        random_gaussian_normal[976] = 16'd126;
        random_gaussian_normal[977] = 16'd1;
        random_gaussian_normal[978] = 16'd45;
        random_gaussian_normal[979] = 16'd378;
        random_gaussian_normal[980] = 16'd35;
        random_gaussian_normal[981] = 16'd31;
        random_gaussian_normal[982] = 16'd179;
        random_gaussian_normal[983] = 16'd62;
        random_gaussian_normal[984] = 16'd236;
        random_gaussian_normal[985] = 16'd166;
        random_gaussian_normal[986] = 16'd42;
        random_gaussian_normal[987] = 16'd481;
        random_gaussian_normal[988] = 16'd140;
        random_gaussian_normal[989] = 16'd247;
        random_gaussian_normal[990] = 16'd132;
        random_gaussian_normal[991] = 16'd253;
        random_gaussian_normal[992] = 16'd314;
        random_gaussian_normal[993] = 16'd398;
        random_gaussian_normal[994] = 16'd8;
        random_gaussian_normal[995] = 16'd35;
        random_gaussian_normal[996] = 16'd540;
        random_gaussian_normal[997] = 16'd31;
        random_gaussian_normal[998] = 16'd5;
        random_gaussian_normal[999] = 16'd232;
        random_gaussian_normal[1000] = 16'd6;
        random_gaussian_normal[1001] = 16'd21;
        random_gaussian_normal[1002] = 16'd123;
        random_gaussian_normal[1003] = 16'd73;
        random_gaussian_normal[1004] = 16'd307;
        random_gaussian_normal[1005] = 16'd114;
        random_gaussian_normal[1006] = 16'd457;
        random_gaussian_normal[1007] = 16'd345;
        random_gaussian_normal[1008] = 16'd223;
        random_gaussian_normal[1009] = 16'd305;
        random_gaussian_normal[1010] = 16'd193;
        random_gaussian_normal[1011] = 16'd179;
        random_gaussian_normal[1012] = 16'd86;
        random_gaussian_normal[1013] = 16'd16;
        random_gaussian_normal[1014] = 16'd67;
        random_gaussian_normal[1015] = 16'd167;
        random_gaussian_normal[1016] = 16'd208;
        random_gaussian_normal[1017] = 16'd194;
        random_gaussian_normal[1018] = 16'd179;
        random_gaussian_normal[1019] = 16'd298;
        random_gaussian_normal[1020] = 16'd175;
        random_gaussian_normal[1021] = 16'd288;
        random_gaussian_normal[1022] = 16'd164;
        random_gaussian_normal[1023] = 16'd203;
    end
    wire signed [15:0] random_gaussian_normal_ori1;
    assign random_gaussian_normal_ori1 = random_gaussian_normal[addr1[9:0]];
    assign random_gaussian_normal_o1 = (random_gaussian_normal_ori1[0] == 1'b1) ? -random_gaussian_normal_ori1[15:1] : random_gaussian_normal_ori1[15:1];

    wire signed [15:0] random_gaussian_normal_ori2;
    assign random_gaussian_normal_ori2 = random_gaussian_normal[addr2[9:0]];
    assign random_gaussian_normal_o2 = (random_gaussian_normal_ori2[0] == 1'b1) ? -random_gaussian_normal_ori2[15:1] : random_gaussian_normal_ori2[15:1];
endmodule